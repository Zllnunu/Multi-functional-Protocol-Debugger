`ifndef DEFINE_VH
`define DEFINE_VH
`define module_name CAN_Top
`define REG
`endif
