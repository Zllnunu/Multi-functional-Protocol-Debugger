`ifndef DEFINE_VH
`define DEFINE_VH
`define module_name CAN_TOP
`define REG
`endif
